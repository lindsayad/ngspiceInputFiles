Alex simple equivalent circuit model of a capacitor
*
* This circuit contains only Berkeley SPICE3 components.
*
* The circuit is an AC coupled transistor amplifier with
* a sinewave input at node "1", a gain of approximately -3.9,
* and output on node "coll".
*
*.tran .005s 2.6673s
.tran 5e0s 5e3s
*
vcc vccTerm 0 10.0
r1 vccTerm r1Term 1MEG 
vdummy0 r1Term vPlas 0.0 
c1 vPlas c1Term 1000uF 
*
s1 vPlas s1Term vPlas 0 smodel1 ON
.MODEL smodel1 SW(VT=5.0 VH=0.0 RON=.9999MEG ROFF=1.0001MEG)
*
vdummy1 c1Term 0 0.0 
vdummy2 s1Term 0 0.0
*
.ic v(vccTerm)=0 v(r1Term)=0 v(vPlas)=0 v(c1Term)=0 v(s1Term)=0
*
*.options TRTOL=100.0 CHGTOL=1.e-16
*
.end


